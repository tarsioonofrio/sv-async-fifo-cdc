module async_fifo
  #(
    parameter BITS=32, // Width of each FIFO entry.
    parameter SIZE=16  // Number of entries. **Recommended: power-of-two** for simpler pointer logic.
  )
  (
    // Write Domain
    input  logic wr_clk,             // Write clock
    input  logic wr_rst_n,           // Active-low write reset (async or sync — see notes)
    input  logic wr_en,              // Write request (one entry per cycle when accepted)
    input  logic [BITS-1:0] wr_data, // Data to write
    output logic wr_full,            // FIFO full flag (do not write when 1)
    // output logic wr_almost_full,          // (Optional) Programmable threshold
    // output logic wr_level,                // (Optional) Approximate fill level (write domain view)
    // Read Domain
    input  logic rd_clk,             // Read clock
    input  logic rd_rst_n,           // Active-low read reset
    input  logic rd_en,              // Read request (one entry per cycle when accepted)
    output logic [BITS-1:0] rd_data, // Data read
    output logic rd_empty            // FIFO empty flag (do not read when 1)
    // output logic rd_almost_empty,         // (Optional) Programmable threshold
    // output logic rd_level,                // (Optional) Approximate fill level (read domain view)
    );


localparam SIZE_LOG2 = $clog2(SIZE);

logic [SIZE-1:0][BITS-1:0] fifo;

logic [SIZE_LOG2:0] wr_ptr_bin;
logic [SIZE_LOG2:0] wr_ptr_bin_next;
logic [SIZE_LOG2:0] wr_ptr_gray;
logic [SIZE_LOG2:0] wr_ptr_bin_sync;
logic [SIZE_LOG2:0] wr_ptr_gray_sync1;
logic [SIZE_LOG2:0] wr_ptr_gray_sync2;

logic [SIZE_LOG2:0] rd_ptr_bin;
logic [SIZE_LOG2:0] rd_ptr_bin_next;
logic [SIZE_LOG2:0] rd_ptr_gray;
logic [SIZE_LOG2:0] rd_ptr_bin_sync;
logic [SIZE_LOG2:0] rd_ptr_gray_sync1;
logic [SIZE_LOG2:0] rd_ptr_gray_sync2;

logic logic_wr_full;
logic logic_rd_empty;


always_ff @(posedge wr_clk) begin
  if (!wr_rst_n) begin
    wr_ptr_bin <= 0;
    wr_ptr_gray <= 0;
  end else if (wr_en && !logic_wr_full) begin
    fifo[wr_ptr_bin[SIZE_LOG2-1:0]] <= wr_data;
    wr_ptr_bin <= wr_ptr_bin + 1;
  end
  wr_ptr_gray <= (wr_ptr_bin_next >> 1) ^ wr_ptr_bin_next;
end
assign wr_ptr_bin_next = wr_ptr_bin + (SIZE_LOG2+1)'(wr_en && !logic_wr_full);

always_ff @(posedge rd_clk) begin
  if (!rd_rst_n) begin
    rd_ptr_bin <= 0;
    rd_ptr_gray <= 0;
  end else if (rd_en && !logic_rd_empty) begin
    rd_data <= fifo[rd_ptr_bin[SIZE_LOG2-1:0]];
    rd_ptr_bin <= rd_ptr_bin + 1;
  end
  rd_ptr_gray <= (rd_ptr_bin_next >> 1) ^ rd_ptr_bin_next;
end
assign rd_ptr_bin_next = rd_ptr_bin + (SIZE_LOG2+1)'(rd_en && !logic_rd_empty);


always_ff @(posedge wr_clk) begin
  if (!wr_rst_n) begin
    rd_ptr_gray_sync1 <= 0;
    rd_ptr_gray_sync2 <= 0;
  end else begin
    rd_ptr_gray_sync1 <= rd_ptr_gray;
    rd_ptr_gray_sync2 <= rd_ptr_gray_sync1;
  end
end

always_ff @(posedge rd_clk) begin
  if (!rd_rst_n) begin
    wr_ptr_gray_sync1 <= 0;
    wr_ptr_gray_sync2 <= 0;
  end else begin
    wr_ptr_gray_sync1 <= wr_ptr_gray;
    wr_ptr_gray_sync2 <= wr_ptr_gray_sync1;
  end
end

generate
  for (genvar i = 0; i < SIZE_LOG2+1; i++) begin: gen_wr_ptr_bin_sync
    assign wr_ptr_bin_sync[i] = ^(wr_ptr_gray_sync2 >> i);
  end

  for (genvar i = 0; i < SIZE_LOG2+1; i++) begin: gen_rd_ptr_bin_sync
    assign rd_ptr_bin_sync[i] = ^(rd_ptr_gray_sync2 >> i);
  end
endgenerate

assign logic_rd_empty = wr_ptr_bin_sync[SIZE_LOG2:0] == rd_ptr_bin[SIZE_LOG2:0];
assign rd_empty = logic_rd_empty;

assign logic_wr_full = (wr_ptr_bin[SIZE_LOG2] != rd_ptr_bin_sync[SIZE_LOG2]) && (wr_ptr_bin[SIZE_LOG2-1:0] == rd_ptr_bin_sync[SIZE_LOG2-1:0]);
assign wr_full = logic_wr_full;

endmodule
